module tb;
input a,b;
output q;
asign q=a|b;
;

