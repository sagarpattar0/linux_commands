rfoufuug
